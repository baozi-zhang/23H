//&----------------------------------------------------------------------------------------
//& 模块名: DA_APMPLITUDE
//& 文件名: DA_APMPLITUDE.v
//& 作  者: 左岚
//& 日  期: 2025-07-18
//&
//& 功  能: DA输出幅度设定模块。该模块提供两个写寄存器，用于通过总线设置两路
//&         DAC（数模转换器）的12位输出幅度值。
//&
//& 设计说明:
//& 1. **重要警告**: 此代码在组合逻辑块(always @(*))中使用了非阻塞赋值(<=)。
//&    这会综合成锁存器(Latch)，而不是推荐使用的时钟同步寄存器(Flip-Flop)。
//&    锁存器对输入毛刺敏感，可能导致不可预测的行为和时序收敛困难。
//&    标准的寄存器设计应在时钟沿触发的 `always` 块中实现。
//& 2. 此模块使用了非标准的双数据总线接口(DATA_ina, DATA_inb)。
//&----------------------------------------------------------------------------------------

module DA_APMPLITUDE #(
    // --- 参数定义 (地址映射) ---
    parameter ADDR14 = 16'h000E,  // DA通道1 幅度值写入地址
    parameter ADDR15 = 16'h000F   // DA通道2 幅度值写入地址
) (
    // --- 端口定义 ---
    // -- 总线控制信号
    input             CS,        // 片选信号，低电平有效
    input             WR_EN,     // 写使能信号，高电平有效
    // -- 数据输入 (非标准接口)
    input      [15:0] DATA_ina,  // 对应地址ADDR14的16位数据输入
    input      [15:0] DATA_inb,  // 对应地址ADDR15的16位数据输入
    // -- 总线地址输入
    input      [15:0] ADDR,      // 16位地址总线
    // -- 寄存器输出 (将作为锁存器实现)
    output reg [11:0] DA1_OUTA,  // DA通道1的12位幅度输出值
    output reg [11:0] DA2_OUTB   // DA通道2的12位幅度输出值
);

  // --- 逻辑实现 ---
  // **警告**: 这是一个组合逻辑块，但使用了非阻塞赋值(<=)，会综合成锁存器。
  always @(*) begin
    // 当片选有效(CS为低)且写使能有效(WR_EN为高)时，执行写操作
    if (!CS && WR_EN) begin
      // 根据地址ADDR，将对应数据总线的低12位锁存到输出寄存器中
      case (ADDR)
        // 地址为ADDR14时，锁存DATA_ina的低12位到DA1_OUTA
        ADDR14: DA1_OUTA <= DATA_ina[11:0];
        // 地址为ADDR15时，锁存DATA_inb的低12位到DA2_OUTB
        ADDR15: DA2_OUTB <= DATA_inb[11:0];
      endcase
    end
  end

endmodule
