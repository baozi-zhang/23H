//&----------------------------------------------------------------------------------------
//& 模块名: DA_CLK_CTRL
//& 文件名: DA_CLK_CTRL.v
//& 作  者: 左岚
//& 日  期: 2025-07-18
//&
//& 功  能: DA时钟控制模块。该模块实现了两个独立的32位数字控制振荡器 (NCO)，
//&         用于根据输入的32位频率控制字生成指定频率的方波信号。
//&         NCO核心原理: F_out = (F_clk * FREQ_WORD) / 2^32
//&
//& 设计说明:
//& 模块B的最终输出 FREQ_OUT_B_FINAL 具有特殊的逻辑：当两个通道的累加器
//& (ACC_A 和 ACC_B) 的值恰好相等时，输出A通道的信号，否则输出B通道自身的信号。
//& 这种设计可能用于特定的同步或锁相应用，但需注意可能引入的瞬时行为。
//&----------------------------------------------------------------------------------------

module DA_CLK_CTRL (
    // --- 端口定义 ---
    input              CLK,               // 系统主时钟
    input              EN,                // 两个NCO的全局使能信号，高电平有效
    // -- 通道A频率控制字输入
    input       [15:0] FREQAH_W,          // 通道A频率控制字的高16位
    input       [15:0] FREQAL_W,          // 通道A频率控制字的低16位
    // -- 通道B频率控制字输入
    input       [15:0] FREQBH_W,          // 通道B频率控制字的高16位
    input       [15:0] FREQBL_W,          // 通道B频率控制字的低16位
    // -- 频率输出
    output wire        FREQ_OUT_A_FINAL,  // 通道A的最终频率输出
    output wire        FREQ_OUT_B_FINAL   // 通道B的最终频率输出
);

  //----------------------------------------------------------------------------------
  //--                             通道A NCO实现
  //----------------------------------------------------------------------------------
  reg [31:0] FREQ_WORD_A;  // 通道A的32位频率控制字寄存器
  reg [31:0] ACC_A = 32'd0;  // 通道A的32位相位累加器，初始值为0
  reg        FREQ_OUT_A;  // 通道A的原始输出（累加器的最高位）

  // 通道A的相位累加器和输出逻辑
  always @(posedge CLK) begin
    if (EN) begin
      // 当使能有效时，累加器在每个时钟周期增加一个频率控制字的值
      ACC_A <= ACC_A + FREQ_WORD_A;
    end
    // 将累加器的最高位(MSB)作为方波输出。当累加器溢出时，该位会翻转。
    FREQ_OUT_A <= ACC_A[31];
  end

  // 通道A的频率控制字输入寄存器
  // 将输入的16位高低字拼接成一个32位的频率字，并在时钟沿锁存，以确保同步
  always @(posedge CLK) begin
    FREQ_WORD_A <= {FREQAH_W, FREQAL_W};
  end

  //----------------------------------------------------------------------------------
  //--                             通道B NCO实现
  //----------------------------------------------------------------------------------
  reg [31:0] FREQ_WORD_B;  // 通道B的32位频率控制字寄存器
  reg [31:0] ACC_B = 32'd0;  // 通道B的32位相位累加器，初始值为0
  reg        FREQ_OUT_B;  // 通道B的原始输出（累加器的最高位）

  // 通道B的相位累加器和输出逻辑
  always @(posedge CLK) begin
    if (EN) begin
      ACC_B <= ACC_B + FREQ_WORD_B;
    end
    FREQ_OUT_B <= ACC_B[31];
  end

  // 通道B的频率控制字输入寄存器
  always @(posedge CLK) begin
    FREQ_WORD_B <= {FREQBH_W, FREQBL_W};
  end

  //----------------------------------------------------------------------------------
  //--                             最终输出逻辑
  //----------------------------------------------------------------------------------
  // 通道B的最终输出逻辑：当两个累加器值相等时，输出A的信号，否则输出B的信号
  assign FREQ_OUT_B_FINAL = (ACC_B == ACC_A) ? FREQ_OUT_A : FREQ_OUT_B;
  // 通道A的最终输出逻辑：直接输出通道A的原始信号
  assign FREQ_OUT_A_FINAL = FREQ_OUT_A;

endmodule
