//&----------------------------------------------------------------------------------------
//& 模块名: DA_FREQ_WORD
//& 文件名: DA_FREQ_WORD.v
//& 作  者: 左岚
//& 日  期: 2025-07-18
//&
//& 功  能: DA频率字设定模块。该模块包含4个16位的写操作寄存器，用于接收外部总线
//&         写入的频率控制字的高低位。
//&
//& 设计说明:
//& 1. **重要警告**: 此代码在组合逻辑块(always @(*))中使用了非阻塞赋值(<=)。
//&    这会导致综合工具生成锁存器(Latch)，而不是推荐使用的时钟同步寄存器(Flip-Flop)。
//&    锁存器对信号毛刺敏感，在设计中应谨慎使用，因为它可能导致时序问题。
//&    正确的寄存器实现方式应使用时序逻辑块 (例如: always @(posedge clk))。
//& 2. 本模块使用了非标准的总线接口，有四个独立的数据输入端(DATA0-DATA3)。
//&----------------------------------------------------------------------------------------

module DA_FREQ_WORD #(
    // --- 参数定义 (地址映射) ---
    parameter ADDR2 = 16'h0002,  // DA通道1 频率字高16位 写入地址
    parameter ADDR3 = 16'h0003,  // DA通道1 频率字低16位 写入地址
    parameter ADDR4 = 16'h0004,  // DA通道2 频率字高16位 写入地址
    parameter ADDR5 = 16'h0005   // DA通道2 频率字低16位 写入地址
) (
    // --- 端口定义 ---
    // -- 总线控制信号
    input             CS,        // 片选信号，低电平有效
    input             WR_EN,     // 写使能信号，高电平有效
    // -- 数据输入 (非标准接口)
    input      [15:0] DATA0,     // 对应地址ADDR2的数据输入
    input      [15:0] DATA1,     // 对应地址ADDR3的数据输入
    input      [15:0] DATA2,     // 对应地址ADDR4的数据输入
    input      [15:0] DATA3,     // 对应地址ADDR5的数据输入
    // -- 总线地址输入
    input      [15:0] ADDR,      // 16位地址总线
    // -- 寄存器输出 (将作为锁存器实现)
    output reg [15:0] DA1_OUTH,  // 存储DA1频率字的高16位
    output reg [15:0] DA1_OUTL,  // 存储DA1频率字的低16位
    output reg [15:0] DA2_OUTH,  // 存储DA2频率字的高16位
    output reg [15:0] DA2_OUTL   // 存储DA2频率字的低16位
);

  // --- 逻辑实现 ---
  // **警告**: 这是一个组合逻辑块，但使用了非阻塞赋值(<=)，会综合成锁存器。
  always @(*) begin
    // 当片选有效(CS为低)且写使能有效(WR_EN为高)时，执行写操作
    if (!CS && WR_EN) begin
      // 根据地址ADDR，将对应的数据输入锁存到输出寄存器中
      case (ADDR)
        ADDR2: DA1_OUTH <= DATA0;  // 地址为ADDR2时，锁存DATA0
        ADDR3: DA1_OUTL <= DATA1;  // 地址为ADDR3时，锁存DATA1
        ADDR4: DA2_OUTH <= DATA2;  // 地址为ADDR4时，锁存DATA2
        ADDR5: DA2_OUTL <= DATA3;  // 地址为ADDR5时，锁存DATA3
      endcase
    end
  end

endmodule
